// Need to figure out how to use hte memory / store the calculaitons